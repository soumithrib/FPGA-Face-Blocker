// nios_system.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module nios_system (
		inout  wire        I2C_SDAT_to_and_from_the_AV_Config,              //        AV_Config_external_interface.SDAT
		output wire        I2C_SCLK_from_the_AV_Config,                     //                                    .SCLK
		inout  wire [15:0] SRAM_DQ_to_and_from_the_Pixel_Buffer,            //     Pixel_Buffer_external_interface.DQ
		output wire [19:0] SRAM_ADDR_from_the_Pixel_Buffer,                 //                                    .ADDR
		output wire        SRAM_LB_N_from_the_Pixel_Buffer,                 //                                    .LB_N
		output wire        SRAM_UB_N_from_the_Pixel_Buffer,                 //                                    .UB_N
		output wire        SRAM_CE_N_from_the_Pixel_Buffer,                 //                                    .CE_N
		output wire        SRAM_OE_N_from_the_Pixel_Buffer,                 //                                    .OE_N
		output wire        SRAM_WE_N_from_the_Pixel_Buffer,                 //                                    .WE_N
		output wire        VGA_CLK_from_the_VGA_Controller,                 //   VGA_Controller_external_interface.CLK
		output wire        VGA_HS_from_the_VGA_Controller,                  //                                    .HS
		output wire        VGA_VS_from_the_VGA_Controller,                  //                                    .VS
		output wire        VGA_BLANK_from_the_VGA_Controller,               //                                    .BLANK
		output wire        VGA_SYNC_from_the_VGA_Controller,                //                                    .SYNC
		output wire [7:0]  VGA_R_from_the_VGA_Controller,                   //                                    .R
		output wire [7:0]  VGA_G_from_the_VGA_Controller,                   //                                    .G
		output wire [7:0]  VGA_B_from_the_VGA_Controller,                   //                                    .B
		input  wire        TD_CLK27_to_the_Video_In_Decoder,                // Video_In_Decoder_external_interface.TD_CLK27
		input  wire [7:0]  TD_DATA_to_the_Video_In_Decoder,                 //                                    .TD_DATA
		input  wire        TD_HS_to_the_Video_In_Decoder,                   //                                    .TD_HS
		input  wire        TD_VS_to_the_Video_In_Decoder,                   //                                    .TD_VS
		input  wire        Video_In_Decoder_external_interface_clk27_reset, //                                    .clk27_reset
		output wire        TD_RESET_from_the_Video_In_Decoder,              //                                    .TD_RESET
		output wire        overflow_flag_from_the_Video_In_Decoder,         //                                    .overflow_flag
		input  wire        clk_clk,                                         //                                 clk.clk
		input  wire [1:0]  pixel_processor_dma_key_n,                       //                 pixel_processor_dma.key_n
		input  wire [17:0] pixel_processor_dma_switch,                      //                                    .switch
		input  wire        reset_reset_n                                    //                               reset.reset_n
	);

	wire         chroma_resampler_avalon_chroma_source_valid;                        // Chroma_Resampler:stream_out_valid -> Color_Space_Converter:stream_in_valid
	wire  [23:0] chroma_resampler_avalon_chroma_source_data;                         // Chroma_Resampler:stream_out_data -> Color_Space_Converter:stream_in_data
	wire         chroma_resampler_avalon_chroma_source_ready;                        // Color_Space_Converter:stream_in_ready -> Chroma_Resampler:stream_out_ready
	wire         chroma_resampler_avalon_chroma_source_startofpacket;                // Chroma_Resampler:stream_out_startofpacket -> Color_Space_Converter:stream_in_startofpacket
	wire         chroma_resampler_avalon_chroma_source_endofpacket;                  // Chroma_Resampler:stream_out_endofpacket -> Color_Space_Converter:stream_in_endofpacket
	wire         video_clipper_avalon_clipper_source_valid;                          // Video_Clipper:stream_out_valid -> Video_Scaler:stream_in_valid
	wire  [15:0] video_clipper_avalon_clipper_source_data;                           // Video_Clipper:stream_out_data -> Video_Scaler:stream_in_data
	wire         video_clipper_avalon_clipper_source_ready;                          // Video_Scaler:stream_in_ready -> Video_Clipper:stream_out_ready
	wire         video_clipper_avalon_clipper_source_startofpacket;                  // Video_Clipper:stream_out_startofpacket -> Video_Scaler:stream_in_startofpacket
	wire         video_clipper_avalon_clipper_source_endofpacket;                    // Video_Clipper:stream_out_endofpacket -> Video_Scaler:stream_in_endofpacket
	wire         color_space_converter_avalon_csc_source_valid;                      // Color_Space_Converter:stream_out_valid -> Video_RGB_Resampler:stream_in_valid
	wire  [23:0] color_space_converter_avalon_csc_source_data;                       // Color_Space_Converter:stream_out_data -> Video_RGB_Resampler:stream_in_data
	wire         color_space_converter_avalon_csc_source_ready;                      // Video_RGB_Resampler:stream_in_ready -> Color_Space_Converter:stream_out_ready
	wire         color_space_converter_avalon_csc_source_startofpacket;              // Color_Space_Converter:stream_out_startofpacket -> Video_RGB_Resampler:stream_in_startofpacket
	wire         color_space_converter_avalon_csc_source_endofpacket;                // Color_Space_Converter:stream_out_endofpacket -> Video_RGB_Resampler:stream_in_endofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_valid;                      // Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire  [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                       // Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire         dual_clock_fifo_avalon_dc_buffer_source_ready;                      // VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	wire         dual_clock_fifo_avalon_dc_buffer_source_startofpacket;              // Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                // Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire         video_in_decoder_avalon_decoder_source_valid;                       // Video_In_Decoder:stream_out_valid -> Chroma_Resampler:stream_in_valid
	wire  [15:0] video_in_decoder_avalon_decoder_source_data;                        // Video_In_Decoder:stream_out_data -> Chroma_Resampler:stream_in_data
	wire         video_in_decoder_avalon_decoder_source_ready;                       // Chroma_Resampler:stream_in_ready -> Video_In_Decoder:stream_out_ready
	wire         video_in_decoder_avalon_decoder_source_startofpacket;               // Video_In_Decoder:stream_out_startofpacket -> Chroma_Resampler:stream_in_startofpacket
	wire         video_in_decoder_avalon_decoder_source_endofpacket;                 // Video_In_Decoder:stream_out_endofpacket -> Chroma_Resampler:stream_in_endofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_valid;                         // Pixel_Buffer_DMA:stream_valid -> Pixel_RGB_Resampler:stream_in_valid
	wire  [15:0] pixel_buffer_dma_avalon_pixel_source_data;                          // Pixel_Buffer_DMA:stream_data -> Pixel_RGB_Resampler:stream_in_data
	wire         pixel_buffer_dma_avalon_pixel_source_ready;                         // Pixel_RGB_Resampler:stream_in_ready -> Pixel_Buffer_DMA:stream_ready
	wire         pixel_buffer_dma_avalon_pixel_source_startofpacket;                 // Pixel_Buffer_DMA:stream_startofpacket -> Pixel_RGB_Resampler:stream_in_startofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_endofpacket;                   // Pixel_Buffer_DMA:stream_endofpacket -> Pixel_RGB_Resampler:stream_in_endofpacket
	wire         video_rgb_resampler_avalon_rgb_source_valid;                        // Video_RGB_Resampler:stream_out_valid -> Video_Clipper:stream_in_valid
	wire  [15:0] video_rgb_resampler_avalon_rgb_source_data;                         // Video_RGB_Resampler:stream_out_data -> Video_Clipper:stream_in_data
	wire         video_rgb_resampler_avalon_rgb_source_ready;                        // Video_Clipper:stream_in_ready -> Video_RGB_Resampler:stream_out_ready
	wire         video_rgb_resampler_avalon_rgb_source_startofpacket;                // Video_RGB_Resampler:stream_out_startofpacket -> Video_Clipper:stream_in_startofpacket
	wire         video_rgb_resampler_avalon_rgb_source_endofpacket;                  // Video_RGB_Resampler:stream_out_endofpacket -> Video_Clipper:stream_in_endofpacket
	wire         pixel_rgb_resampler_avalon_rgb_source_valid;                        // Pixel_RGB_Resampler:stream_out_valid -> Pixel_Scaler:stream_in_valid
	wire  [29:0] pixel_rgb_resampler_avalon_rgb_source_data;                         // Pixel_RGB_Resampler:stream_out_data -> Pixel_Scaler:stream_in_data
	wire         pixel_rgb_resampler_avalon_rgb_source_ready;                        // Pixel_Scaler:stream_in_ready -> Pixel_RGB_Resampler:stream_out_ready
	wire         pixel_rgb_resampler_avalon_rgb_source_startofpacket;                // Pixel_RGB_Resampler:stream_out_startofpacket -> Pixel_Scaler:stream_in_startofpacket
	wire         pixel_rgb_resampler_avalon_rgb_source_endofpacket;                  // Pixel_RGB_Resampler:stream_out_endofpacket -> Pixel_Scaler:stream_in_endofpacket
	wire         pixel_scaler_avalon_scaler_source_valid;                            // Pixel_Scaler:stream_out_valid -> Dual_Clock_FIFO:stream_in_valid
	wire  [29:0] pixel_scaler_avalon_scaler_source_data;                             // Pixel_Scaler:stream_out_data -> Dual_Clock_FIFO:stream_in_data
	wire         pixel_scaler_avalon_scaler_source_ready;                            // Dual_Clock_FIFO:stream_in_ready -> Pixel_Scaler:stream_out_ready
	wire         pixel_scaler_avalon_scaler_source_startofpacket;                    // Pixel_Scaler:stream_out_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	wire         pixel_scaler_avalon_scaler_source_endofpacket;                      // Pixel_Scaler:stream_out_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	wire         video_scaler_avalon_scaler_source_valid;                            // Video_Scaler:stream_out_valid -> Pixel_Processor_DMA:stream_valid
	wire  [15:0] video_scaler_avalon_scaler_source_data;                             // Video_Scaler:stream_out_data -> Pixel_Processor_DMA:stream_data
	wire         video_scaler_avalon_scaler_source_ready;                            // Pixel_Processor_DMA:stream_ready -> Video_Scaler:stream_out_ready
	wire         video_scaler_avalon_scaler_source_startofpacket;                    // Video_Scaler:stream_out_startofpacket -> Pixel_Processor_DMA:stream_startofpacket
	wire         video_scaler_avalon_scaler_source_endofpacket;                      // Video_Scaler:stream_out_endofpacket -> Pixel_Processor_DMA:stream_endofpacket
	wire         video_pll_0_vga_clk_clk;                                            // video_pll_0:vga_clk_clk -> [Dual_Clock_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_002:clk]
	wire         pixel_processor_dma_avalon_master_waitrequest;                      // mm_interconnect_0:Pixel_Processor_DMA_avalon_master_waitrequest -> Pixel_Processor_DMA:master_waitrequest
	wire  [31:0] pixel_processor_dma_avalon_master_address;                          // Pixel_Processor_DMA:master_address -> mm_interconnect_0:Pixel_Processor_DMA_avalon_master_address
	wire         pixel_processor_dma_avalon_master_write;                            // Pixel_Processor_DMA:master_write -> mm_interconnect_0:Pixel_Processor_DMA_avalon_master_write
	wire  [15:0] pixel_processor_dma_avalon_master_writedata;                        // Pixel_Processor_DMA:master_writedata -> mm_interconnect_0:Pixel_Processor_DMA_avalon_master_writedata
	wire         pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;               // mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_waitrequest -> Pixel_Buffer_DMA:master_waitrequest
	wire  [15:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                  // mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_readdata -> Pixel_Buffer_DMA:master_readdata
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                   // Pixel_Buffer_DMA:master_address -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_address
	wire         pixel_buffer_dma_avalon_pixel_dma_master_read;                      // Pixel_Buffer_DMA:master_read -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_read
	wire         pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;             // mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_readdatavalid -> Pixel_Buffer_DMA:master_readdatavalid
	wire         pixel_buffer_dma_avalon_pixel_dma_master_lock;                      // Pixel_Buffer_DMA:master_arbiterlock -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_lock
	wire  [31:0] cpu_data_master_readdata;                                           // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                                        // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                                        // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [21:0] cpu_data_master_address;                                            // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                         // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                               // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                              // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                          // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                    // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                                 // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [21:0] cpu_instruction_master_address;                                     // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                        // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata;          // Pixel_Buffer:readdata -> mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_address;           // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_address -> Pixel_Buffer:address
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_read;              // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_read -> Pixel_Buffer:read
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable;        // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_byteenable -> Pixel_Buffer:byteenable
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid;     // Pixel_Buffer:readdatavalid -> mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_write;             // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_write -> Pixel_Buffer:write
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata;         // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_writedata -> Pixel_Buffer:writedata
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_readdata;        // AV_Config:readdata -> mm_interconnect_0:AV_Config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest;     // AV_Config:waitrequest -> mm_interconnect_0:AV_Config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_av_config_avalon_av_config_slave_address;         // mm_interconnect_0:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_read;            // mm_interconnect_0:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	wire   [3:0] mm_interconnect_0_av_config_avalon_av_config_slave_byteenable;      // mm_interconnect_0:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_write;           // mm_interconnect_0:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_writedata;       // mm_interconnect_0:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata;   // Pixel_Buffer_DMA:slave_readdata -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address;    // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_address -> Pixel_Buffer_DMA:slave_address
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read;       // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_read -> Pixel_Buffer_DMA:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable; // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_byteenable -> Pixel_Buffer_DMA:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write;      // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_write -> Pixel_Buffer_DMA:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata;  // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_writedata -> Pixel_Buffer_DMA:slave_writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                   // CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                // CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                // mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                    // mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                       // mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                 // mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                      // mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                  // mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                      // mm_interconnect_0:Onchip_Memory_s1_chipselect -> Onchip_Memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                        // Onchip_Memory:readdata -> mm_interconnect_0:Onchip_Memory_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory_s1_address;                         // mm_interconnect_0:Onchip_Memory_s1_address -> Onchip_Memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                      // mm_interconnect_0:Onchip_Memory_s1_byteenable -> Onchip_Memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                           // mm_interconnect_0:Onchip_Memory_s1_write -> Onchip_Memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                       // mm_interconnect_0:Onchip_Memory_s1_writedata -> Onchip_Memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                           // mm_interconnect_0:Onchip_Memory_s1_clken -> Onchip_Memory:clken
	wire  [31:0] cpu_d_irq_irq;                                                      // irq_mapper:sender_irq -> CPU:d_irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [AV_Config:reset, Chroma_Resampler:reset, Color_Space_Converter:reset, Dual_Clock_FIFO:reset_stream_in, Pixel_Buffer:reset, Pixel_Buffer_DMA:reset, Pixel_Processor_DMA:reset, Pixel_RGB_Resampler:reset, Pixel_Scaler:reset, Video_Clipper:reset, Video_In_Decoder:reset, Video_RGB_Resampler:reset, Video_Scaler:reset, mm_interconnect_0:Pixel_Processor_DMA_reset_reset_bridge_in_reset_reset, video_pll_0:ref_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [CPU:reset_n, Onchip_Memory:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [CPU:reset_req, Onchip_Memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                  // CPU:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [Dual_Clock_FIFO:reset_stream_out, VGA_Controller:reset]
	wire         video_pll_0_reset_source_reset;                                     // video_pll_0:reset_source_reset -> rst_controller_002:reset_in0

	nios_system_AV_Config av_config (
		.clk         (clk_clk),                                                        //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //                  reset.reset
		.address     (mm_interconnect_0_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (I2C_SDAT_to_and_from_the_AV_Config),                             //     external_interface.export
		.I2C_SCLK    (I2C_SCLK_from_the_AV_Config)                                     //                       .export
	);

	nios_system_CPU cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	nios_system_Chroma_Resampler chroma_resampler (
		.clk                      (clk_clk),                                              //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                       //                reset.reset
		.stream_in_startofpacket  (video_in_decoder_avalon_decoder_source_startofpacket), //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (video_in_decoder_avalon_decoder_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_in_decoder_avalon_decoder_source_valid),         //                     .valid
		.stream_in_ready          (video_in_decoder_avalon_decoder_source_ready),         //                     .ready
		.stream_in_data           (video_in_decoder_avalon_decoder_source_data),          //                     .data
		.stream_out_ready         (chroma_resampler_avalon_chroma_source_ready),          // avalon_chroma_source.ready
		.stream_out_startofpacket (chroma_resampler_avalon_chroma_source_startofpacket),  //                     .startofpacket
		.stream_out_endofpacket   (chroma_resampler_avalon_chroma_source_endofpacket),    //                     .endofpacket
		.stream_out_valid         (chroma_resampler_avalon_chroma_source_valid),          //                     .valid
		.stream_out_data          (chroma_resampler_avalon_chroma_source_data)            //                     .data
	);

	nios_system_Color_Space_Converter color_space_converter (
		.clk                      (clk_clk),                                               //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //             reset.reset
		.stream_in_startofpacket  (chroma_resampler_avalon_chroma_source_startofpacket),   //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (chroma_resampler_avalon_chroma_source_endofpacket),     //                  .endofpacket
		.stream_in_valid          (chroma_resampler_avalon_chroma_source_valid),           //                  .valid
		.stream_in_ready          (chroma_resampler_avalon_chroma_source_ready),           //                  .ready
		.stream_in_data           (chroma_resampler_avalon_chroma_source_data),            //                  .data
		.stream_out_ready         (color_space_converter_avalon_csc_source_ready),         // avalon_csc_source.ready
		.stream_out_startofpacket (color_space_converter_avalon_csc_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (color_space_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (color_space_converter_avalon_csc_source_valid),         //                  .valid
		.stream_out_data          (color_space_converter_avalon_csc_source_data)           //                  .data
	);

	nios_system_Dual_Clock_FIFO dual_clock_fifo (
		.clk_stream_in            (clk_clk),                                               //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                        //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                               //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                    //        reset_stream_out.reset
		.stream_in_ready          (pixel_scaler_avalon_scaler_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (pixel_scaler_avalon_scaler_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (pixel_scaler_avalon_scaler_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (pixel_scaler_avalon_scaler_source_valid),               //                        .valid
		.stream_in_data           (pixel_scaler_avalon_scaler_source_data),                //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_Onchip_Memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)         //       .reset_req
	);

	nios_system_Pixel_Buffer pixel_buffer (
		.clk           (clk_clk),                                                        //                clk.clk
		.reset         (rst_controller_reset_out_reset),                                 //              reset.reset
		.SRAM_DQ       (SRAM_DQ_to_and_from_the_Pixel_Buffer),                           // external_interface.export
		.SRAM_ADDR     (SRAM_ADDR_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_LB_N     (SRAM_LB_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_UB_N     (SRAM_UB_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_CE_N     (SRAM_CE_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_OE_N     (SRAM_OE_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_WE_N     (SRAM_WE_N_from_the_Pixel_Buffer),                                //                   .export
		.address       (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_Pixel_Buffer_DMA pixel_buffer_dma (
		.clk                  (clk_clk),                                                            //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                     //                   reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                           //                        .data
	);

	pixel_processor_DMA pixel_processor_dma (
		.clk                  (clk_clk),                                         //                 clock.clk
		.reset                (rst_controller_reset_out_reset),                  //                 reset.reset
		.slave_address        (),                                                //                 slave.address
		.slave_byteenable     (),                                                //                      .byteenable
		.slave_read           (),                                                //                      .read
		.slave_write          (),                                                //                      .write
		.slave_writedata      (),                                                //                      .writedata
		.slave_readdata       (),                                                //                      .readdata
		.stream_data          (video_scaler_avalon_scaler_source_data),          // avalon_streaming_sink.data
		.stream_endofpacket   (video_scaler_avalon_scaler_source_endofpacket),   //                      .endofpacket
		.stream_ready         (video_scaler_avalon_scaler_source_ready),         //                      .ready
		.stream_startofpacket (video_scaler_avalon_scaler_source_startofpacket), //                      .startofpacket
		.stream_valid         (video_scaler_avalon_scaler_source_valid),         //                      .valid
		.master_waitrequest   (pixel_processor_dma_avalon_master_waitrequest),   //         avalon_master.waitrequest
		.master_address       (pixel_processor_dma_avalon_master_address),       //                      .address
		.master_write         (pixel_processor_dma_avalon_master_write),         //                      .write
		.master_writedata     (pixel_processor_dma_avalon_master_writedata),     //                      .writedata
		.key_n                (pixel_processor_dma_key_n),                       //           conduit_end.key_n
		.s                    (pixel_processor_dma_switch)                       //                      .switch
	);

	nios_system_Pixel_RGB_Resampler pixel_rgb_resampler (
		.clk                      (clk_clk),                                             //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket),  //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),    //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),          //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),          //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),           //                  .data
		.stream_out_ready         (pixel_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (pixel_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (pixel_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (pixel_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios_system_Pixel_Scaler pixel_scaler (
		.clk                      (clk_clk),                                             //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                reset.reset
		.stream_in_startofpacket  (pixel_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (pixel_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (pixel_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (pixel_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (pixel_scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (pixel_scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (pixel_scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (pixel_scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (pixel_scaler_avalon_scaler_source_data)               //                     .data
	);

	nios_system_VGA_Controller vga_controller (
		.clk           (video_pll_0_vga_clk_clk),                               //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                    //              reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (VGA_CLK_from_the_VGA_Controller),                       // external_interface.export
		.VGA_HS        (VGA_HS_from_the_VGA_Controller),                        //                   .export
		.VGA_VS        (VGA_VS_from_the_VGA_Controller),                        //                   .export
		.VGA_BLANK     (VGA_BLANK_from_the_VGA_Controller),                     //                   .export
		.VGA_SYNC      (VGA_SYNC_from_the_VGA_Controller),                      //                   .export
		.VGA_R         (VGA_R_from_the_VGA_Controller),                         //                   .export
		.VGA_G         (VGA_G_from_the_VGA_Controller),                         //                   .export
		.VGA_B         (VGA_B_from_the_VGA_Controller)                          //                   .export
	);

	nios_system_Video_Clipper video_clipper (
		.clk                      (clk_clk),                                             //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                 reset.reset
		.stream_in_data           (video_rgb_resampler_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_rgb_resampler_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (video_rgb_resampler_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (video_rgb_resampler_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (video_clipper_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (video_clipper_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (video_clipper_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (video_clipper_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (video_clipper_avalon_clipper_source_valid)            //                      .valid
	);

	nios_system_Video_In_Decoder video_in_decoder (
		.clk                      (clk_clk),                                              //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                       //                 reset.reset
		.stream_out_ready         (video_in_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_in_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_in_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_in_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_in_decoder_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (TD_CLK27_to_the_Video_In_Decoder),                     //    external_interface.export
		.TD_DATA                  (TD_DATA_to_the_Video_In_Decoder),                      //                      .export
		.TD_HS                    (TD_HS_to_the_Video_In_Decoder),                        //                      .export
		.TD_VS                    (TD_VS_to_the_Video_In_Decoder),                        //                      .export
		.clk27_reset              (Video_In_Decoder_external_interface_clk27_reset),      //                      .export
		.TD_RESET                 (TD_RESET_from_the_Video_In_Decoder),                   //                      .export
		.overflow_flag            (overflow_flag_from_the_Video_In_Decoder)               //                      .export
	);

	nios_system_Video_RGB_Resampler video_rgb_resampler (
		.clk                      (clk_clk),                                               //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //             reset.reset
		.stream_in_startofpacket  (color_space_converter_avalon_csc_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (color_space_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (color_space_converter_avalon_csc_source_valid),         //                  .valid
		.stream_in_ready          (color_space_converter_avalon_csc_source_ready),         //                  .ready
		.stream_in_data           (color_space_converter_avalon_csc_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_avalon_rgb_source_ready),           // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_avalon_rgb_source_startofpacket),   //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_avalon_rgb_source_endofpacket),     //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_avalon_rgb_source_valid),           //                  .valid
		.stream_out_data          (video_rgb_resampler_avalon_rgb_source_data)             //                  .data
	);

	nios_system_Video_Scaler video_scaler (
		.clk                      (clk_clk),                                           //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                    //                reset.reset
		.stream_in_startofpacket  (video_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_scaler_avalon_scaler_source_data)             //                     .data
	);

	nios_system_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (rst_controller_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)  // reset_source.reset
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                          (clk_clk),                                                            //                                       clk_0_clk.clk
		.CPU_reset_n_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                                 //               CPU_reset_n_reset_bridge_in_reset.reset
		.Pixel_Processor_DMA_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                     // Pixel_Processor_DMA_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                                (cpu_data_master_address),                                            //                                 CPU_data_master.address
		.CPU_data_master_waitrequest                            (cpu_data_master_waitrequest),                                        //                                                .waitrequest
		.CPU_data_master_byteenable                             (cpu_data_master_byteenable),                                         //                                                .byteenable
		.CPU_data_master_read                                   (cpu_data_master_read),                                               //                                                .read
		.CPU_data_master_readdata                               (cpu_data_master_readdata),                                           //                                                .readdata
		.CPU_data_master_write                                  (cpu_data_master_write),                                              //                                                .write
		.CPU_data_master_writedata                              (cpu_data_master_writedata),                                          //                                                .writedata
		.CPU_data_master_debugaccess                            (cpu_data_master_debugaccess),                                        //                                                .debugaccess
		.CPU_instruction_master_address                         (cpu_instruction_master_address),                                     //                          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                     (cpu_instruction_master_waitrequest),                                 //                                                .waitrequest
		.CPU_instruction_master_read                            (cpu_instruction_master_read),                                        //                                                .read
		.CPU_instruction_master_readdata                        (cpu_instruction_master_readdata),                                    //                                                .readdata
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //        Pixel_Buffer_DMA_avalon_pixel_dma_master.address
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                                                .waitrequest
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                                                .read
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                                                .readdata
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             //                                                .readdatavalid
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_lock          (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                                                .lock
		.Pixel_Processor_DMA_avalon_master_address              (pixel_processor_dma_avalon_master_address),                          //               Pixel_Processor_DMA_avalon_master.address
		.Pixel_Processor_DMA_avalon_master_waitrequest          (pixel_processor_dma_avalon_master_waitrequest),                      //                                                .waitrequest
		.Pixel_Processor_DMA_avalon_master_write                (pixel_processor_dma_avalon_master_write),                            //                                                .write
		.Pixel_Processor_DMA_avalon_master_writedata            (pixel_processor_dma_avalon_master_writedata),                        //                                                .writedata
		.AV_Config_avalon_av_config_slave_address               (mm_interconnect_0_av_config_avalon_av_config_slave_address),         //                AV_Config_avalon_av_config_slave.address
		.AV_Config_avalon_av_config_slave_write                 (mm_interconnect_0_av_config_avalon_av_config_slave_write),           //                                                .write
		.AV_Config_avalon_av_config_slave_read                  (mm_interconnect_0_av_config_avalon_av_config_slave_read),            //                                                .read
		.AV_Config_avalon_av_config_slave_readdata              (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),        //                                                .readdata
		.AV_Config_avalon_av_config_slave_writedata             (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),       //                                                .writedata
		.AV_Config_avalon_av_config_slave_byteenable            (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),      //                                                .byteenable
		.AV_Config_avalon_av_config_slave_waitrequest           (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest),     //                                                .waitrequest
		.CPU_jtag_debug_module_address                          (mm_interconnect_0_cpu_jtag_debug_module_address),                    //                           CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                            (mm_interconnect_0_cpu_jtag_debug_module_write),                      //                                                .write
		.CPU_jtag_debug_module_read                             (mm_interconnect_0_cpu_jtag_debug_module_read),                       //                                                .read
		.CPU_jtag_debug_module_readdata                         (mm_interconnect_0_cpu_jtag_debug_module_readdata),                   //                                                .readdata
		.CPU_jtag_debug_module_writedata                        (mm_interconnect_0_cpu_jtag_debug_module_writedata),                  //                                                .writedata
		.CPU_jtag_debug_module_byteenable                       (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                 //                                                .byteenable
		.CPU_jtag_debug_module_waitrequest                      (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                //                                                .waitrequest
		.CPU_jtag_debug_module_debugaccess                      (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                //                                                .debugaccess
		.Onchip_Memory_s1_address                               (mm_interconnect_0_onchip_memory_s1_address),                         //                                Onchip_Memory_s1.address
		.Onchip_Memory_s1_write                                 (mm_interconnect_0_onchip_memory_s1_write),                           //                                                .write
		.Onchip_Memory_s1_readdata                              (mm_interconnect_0_onchip_memory_s1_readdata),                        //                                                .readdata
		.Onchip_Memory_s1_writedata                             (mm_interconnect_0_onchip_memory_s1_writedata),                       //                                                .writedata
		.Onchip_Memory_s1_byteenable                            (mm_interconnect_0_onchip_memory_s1_byteenable),                      //                                                .byteenable
		.Onchip_Memory_s1_chipselect                            (mm_interconnect_0_onchip_memory_s1_chipselect),                      //                                                .chipselect
		.Onchip_Memory_s1_clken                                 (mm_interconnect_0_onchip_memory_s1_clken),                           //                                                .clken
		.Pixel_Buffer_avalon_sram_slave_address                 (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),           //                  Pixel_Buffer_avalon_sram_slave.address
		.Pixel_Buffer_avalon_sram_slave_write                   (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),             //                                                .write
		.Pixel_Buffer_avalon_sram_slave_read                    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),              //                                                .read
		.Pixel_Buffer_avalon_sram_slave_readdata                (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),          //                                                .readdata
		.Pixel_Buffer_avalon_sram_slave_writedata               (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),         //                                                .writedata
		.Pixel_Buffer_avalon_sram_slave_byteenable              (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),        //                                                .byteenable
		.Pixel_Buffer_avalon_sram_slave_readdatavalid           (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid),     //                                                .readdatavalid
		.Pixel_Buffer_DMA_avalon_control_slave_address          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //           Pixel_Buffer_DMA_avalon_control_slave.address
		.Pixel_Buffer_DMA_avalon_control_slave_write            (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                                                .write
		.Pixel_Buffer_DMA_avalon_control_slave_read             (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                                                .read
		.Pixel_Buffer_DMA_avalon_control_slave_readdata         (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                                                .readdata
		.Pixel_Buffer_DMA_avalon_control_slave_writedata        (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                                                .writedata
		.Pixel_Buffer_DMA_avalon_control_slave_byteenable       (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable)  //                                                .byteenable
	);

	nios_system_irq_mapper irq_mapper (
		.clk        (clk_clk),                            //       clk.clk
		.reset      (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
